-- Generated PORTMAP Stub File: Created by Capture FPGA Flow
-- Matches PCB component pinout with simulation model
-- Created Saturday, May 25, 2024 19:57:16 GTB Daylight Time

